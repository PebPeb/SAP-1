----------------------------------------------
-- program_counter								--
-- 											--
-- Keeps track of the program location						--
-- 								 			--
-- Original Project : SAP-1					--
-- By: Bryce Keen				 			--
-- 06/30/22 								--
----------------------------------------------


library ieee;
use IEEE.STD_LOGIC_1164.all;


entity program_counter is
	port (
		CLK:		in STD_lOGIC;						-- Clock and LB
	);
end;


architecture program_counter_arch of program_counter is	
  
begin

	-- Logic

	
	-- Output Logic
	
	
end program_counter_arch;
